module IR_MEM (pc_ir,ir);
input [31:0] pc_ir;
output reg [31:0]ir;
reg [31:0] IR_MEM [0:1023];

 integer i;
    initial begin
        for(i = 0; i <=1023; i = i + 1) begin
			IR_MEM[i] = 0;
		end
    end
	 
always @(pc_ir)
begin
ir=IR_MEM[pc_ir];
end

initial 
begin

IR_MEM[0]={7'b0000000,5'b00001,5'b00111,3'b000,5'b00111,7'b0110011};// add 
IR_MEM[1]={7'b1111111,5'b00111,5'b00011,3'b001,5'b11111,7'b1100011};


//IR_MEM[1]={7'b0100000,5'b00010,5'b00001,3'b000,5'b00101,7'b0110011};// sub 
//IR_MEM[2]={7'b0000000,5'b00011,5'b00111,3'b000,5'b00001,7'b0110011};// add 

//IR_MEM[0]={7'b0000000,5'b00110,5'b00100,3'b110,5'b00001,7'b0110011};// or r1,r4,r6
//IR_MEM[1]={7'b0100000,5'b00100,5'b00110,3'b111,5'b00010,7'b0110011};// and r2,r6,r4

//IR_MEM[0]={7'b0000000,5'b00111,5'b00100,3'b000,5'b00001,7'b0010011};// addi r1,r4,7
//IR_MEM[1]={7'b0000000,5'b00011,5'b00111,3'b111,5'b00010,7'b0010011};// andi r2,r7,3

//IR_MEM[0]={7'b0000000,5'b00100,5'b00000,3'b000,5'b00001,7'b0100011};// sb r4,01(r0)
//IR_MEM[0]={7'b0000000,5'b00011,5'b00000,3'b010,5'b00010,7'b0100011};// sw r7,02(r0)

//IR_MEM[0]={7'b0000000,5'b00001,5'b00000,3'b001,5'b00110,7'b0000011};// lw r6,1(r0)
//IR_MEM[1]={7'b0000000,5'b00010,5'b00000,3'b000,5'b00111,7'b0000011};// lb r7,2(r0)




/*
IR_MEM[0]={7'b0000000,5'b00111,5'b00000,3'b000,5'b00110,7'b0010011};// addi r6,r0,7
IR_MEM[1]={7'b0000000,5'b00011,5'b00000,3'b000,5'b00111,7'b0010011};// addi r7,r0,3
IR_MEM[2]={7'b0000000,5'b00000,5'b00000,3'b110,5'b00101,7'b0110011};// dummy instruction
IR_MEM[3]={7'b0000000,5'b00000,5'b00000,3'b110,5'b00101,7'b0110011};// dummy instruction
IR_MEM[4]={7'b0000000,5'b00110,5'b00111,3'b000,5'b00001,7'b0110011};// add r1,r6,r7
*/


//IR_MEM[0]={7'b0000000,5'b00100,5'b00000,3'b010,5'b00001,7'b0100011};
//IR_MEM[1]={7'b0000000,5'b00000,5'b00000,3'b000,5'b00001,7'b1101111};
/*
IR_MEM[0]={7'b0000000,5'b01010,5'b00100,3'b000,5'b00011,7'b0010011};// addi 
IR_MEM[1]={7'b0000000,5'b00111,5'b00110,3'b000,5'b00101,7'b0110011};// add
*/
/*
IR_MEM[2]={7'b1111111,5'b10000,5'b00000,3'b000,5'b00011,7'b0010011};// addi r3,ff0(r0)
IR_MEM[3]={7'b0000000,5'b00001,5'b00001,3'b000,5'b00001,7'b0010011};// addi r3,ff0(r0)
IR_MEM[6]={7'b0000000,5'b01111,5'b00000,3'b000,5'b00110,7'b0010011};// addi r2,00f(r0)
IR_MEM[7]={7'b0000000,5'b01011,5'b00000,3'b000,5'b00111,7'b0010011};// addi r2,00f(r0)
*/
//IR_MEM[4]={7'b1111111,5'b00000,5'b00000,3'b000,5'b11101,7'b1100011};// addi r4,f(r0)

//IR_MEM[5]={  7'b0000000,5'b00001,5'b00001,3'b000,5'b00001,7'b0010011};// addi r3,ff0(r0)
//IR_MEM[5]={7'b0000000,5'b00001,5'b00000,3'b010,5'b00001,7'b0100011};// sw r1,05(r0)
//IR_MEM[6]={7'b0000000,5'b00001,5'b00000,3'b010,5'b00010,7'b0100011};// sw r1,05(r0)
//IR_MEM[7]={7'b0000000,5'b00100,5'b00000,3'b010,5'b00011,7'b0100011};// sw
end

endmodule 
	
